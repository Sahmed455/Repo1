module AND2(
	input in1,
	input in2,
	output Out
	);
//	$display("ADD2 Running!!!");
//	$finish;
	assign Out=in1&in2;

endmodule
