module XOR2(
	input in1,
	input in2,
	output Out
);
assign Out=in1^in2;
endmodule
